module mkmac8(CLK,
	      RST,

	      get_values_multiplicand1,
	      get_values_multiplicand2,
	      get_values_addend,
	      EN_get_values,
	      RDY_get_values,

	      mac_result,
	      RDY_mac_result);
  input  CLK;
  input  RST;

  // action method get_values
  input  [7 : 0] get_values_multiplicand1;
  input  [7 : 0] get_values_multiplicand2;
  input  [7 : 0] get_values_addend;
  input  EN_get_values;
  output RDY_get_values;

  // value method mac_result
  output [15 : 0] mac_result;
  output RDY_mac_result;

  // signals for module outputs
  wire [15 : 0] mac_result;
  wire RDY_get_values, RDY_mac_result;

  // register a
  reg [7 : 0] a;
  wire [7 : 0] a$D_IN;
  wire a$EN;

  // register inp_ready
  reg inp_ready;
  wire inp_ready$D_IN, inp_ready$EN;

  // register m1
  reg [7 : 0] m1;
  wire [7 : 0] m1$D_IN;
  wire m1$EN;

  // register m2
  reg [7 : 0] m2;
  wire [7 : 0] m2$D_IN;
  wire m2$EN;

  // register mac_ready
  reg mac_ready;
  wire mac_ready$D_IN, mac_ready$EN;

  // register resmac
  reg [15 : 0] resmac;
  wire [15 : 0] resmac$D_IN;
  wire resmac$EN;

  // rule scheduling signals
  wire CAN_FIRE_RL_mac,
       CAN_FIRE_get_values,
       WILL_FIRE_RL_mac,
       WILL_FIRE_get_values;

  // remaining internal signals
  wire [31 : 0] _0_CONCAT_m1_MUL_0_CONCAT_m2___d6;
  wire [15 : 0] x__h299, y__h298, y__h300;
  wire NOT_get_values_multiplicand1_EQ_m1_1_2_OR_NOT__ETC___d18;

  // action method get_values
  assign RDY_get_values = 1'd1 ;
  assign CAN_FIRE_get_values = 1'd1 ;
  assign WILL_FIRE_get_values = EN_get_values ;

  // value method mac_result
  assign mac_result = resmac ;
  assign RDY_mac_result = mac_ready ;

  // rule RL_mac
  assign CAN_FIRE_RL_mac = 1'd1 ;
  assign WILL_FIRE_RL_mac = 1'd1 ;

  // register a
  assign a$D_IN = get_values_addend ;
  assign a$EN =
	     EN_get_values &&
	     NOT_get_values_multiplicand1_EQ_m1_1_2_OR_NOT__ETC___d18 ;

  // register inp_ready
  assign inp_ready$D_IN =
	     NOT_get_values_multiplicand1_EQ_m1_1_2_OR_NOT__ETC___d18 ;
  assign inp_ready$EN = EN_get_values ;

  // register m1
  assign m1$D_IN = get_values_multiplicand1 ;
  assign m1$EN =
	     EN_get_values &&
	     NOT_get_values_multiplicand1_EQ_m1_1_2_OR_NOT__ETC___d18 ;

  // register m2
  assign m2$D_IN = get_values_multiplicand2 ;
  assign m2$EN =
	     EN_get_values &&
	     NOT_get_values_multiplicand1_EQ_m1_1_2_OR_NOT__ETC___d18 ;

  // register mac_ready
  assign mac_ready$D_IN = inp_ready ;
  assign mac_ready$EN = 1'd1 ;

  // register resmac
  assign resmac$D_IN = _0_CONCAT_m1_MUL_0_CONCAT_m2___d6[15:0] + y__h298 ;
  assign resmac$EN = inp_ready ;

  // remaining internal signals
  assign NOT_get_values_multiplicand1_EQ_m1_1_2_OR_NOT__ETC___d18 =
	     get_values_multiplicand1 != m1 ||
	     get_values_multiplicand2 != m2 ||
	     get_values_addend != a ;
  assign _0_CONCAT_m1_MUL_0_CONCAT_m2___d6 = x__h299 * y__h300 ;
  assign x__h299 = { 8'd0, m1 } ;
  assign y__h298 = { 8'd0, a } ;
  assign y__h300 = { 8'd0, m2 } ;

  // handling of inlined registers

  always@(posedge CLK)
  begin
    if (RST == 1)
      begin
        a <= 8'd0;
	inp_ready <= 1'd0;
	m1 <= 8'd0;
	m2 <= 8'd0;
	mac_ready <= 1'd0;
	resmac <= 16'd0;
      end
    else
      begin
        if (a$EN) a <= a$D_IN;
	if (inp_ready$EN) inp_ready <= inp_ready$D_IN;
	if (m1$EN) m1 <= m1$D_IN;
	if (m2$EN) m2 <= m2$D_IN;
	if (mac_ready$EN) mac_ready <= mac_ready$D_IN;
	if (resmac$EN) resmac <= resmac$D_IN;
      end
  end

  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    a = 8'hAA;
    inp_ready = 1'h0;
    m1 = 8'hAA;
    m2 = 8'hAA;
    mac_ready = 1'h0;
    resmac = 16'hAAAA;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on
endmodule  // mkmac8

