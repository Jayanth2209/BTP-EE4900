module mkMAC(
         input CLK,
	     input RST,

	     input [63:0] m1,
	     input [63:0] m2,
	     input [63:0] a,
	     input [1:0] mode,
	     input EN_get_values,
	     output RDY_get_values,

	     output [127:0] mac_result,
	     output RDY_mac_result);



endmodule